module gradient(input [7:0] window[0:5][0:5], output [7:0] Gx[0:3][0:3], output [7:0] Gy[0:3][0:3]);

endmodule