module window_gen(input[7:0] pixel,output[7:0] window[0:5][0:5]);

endmodule