module rgb_to_grey(input clk, input[7:0] Rpixel,input[7:0] Gpixel,input[7:0] Bpixel, output[7:0] pixel);

    


endmodule