module(input [7:0] Gx[0:3][0:3], input [7:0] Gy[0:3][0:3], output [7:0] R);
endmodule